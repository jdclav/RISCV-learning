module ALU (
    input CLK,        
    input RESET,      
    input ALU,
    input ALUimm,
    input [31:0] rs1,
    input [31:0] rs2,
    input [2:0] funct3,
    input [6:0] funct7,
    output [31:0] ALUresult
);







endmodule